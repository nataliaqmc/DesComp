library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;    -- Biblioteca IEEE para funções aritméticas

entity logicaDisplays is
    port (
		CLK : in std_logic;
    );
end entity;

architecture comportamento of logicaDisplay is

    begin
      		
end architecture;